** Simple BJT Class A Pre-Amplifier
** Template Class A BJT Amplifier
** Author: Nathan Campos <nathanpc@dreamintech.net>


**
** Circuit
**

** First stage.

* Base
C1 input q1b 2.2u
R1 v+ q1b 47k
R2 q1b 0 10k

* Collector
R3 v+ q1c 5k
C2 q1c output 0.1u

* Emitter
R4 q1e 0 1k

* Transistor
Q1 q1c q1b q1e q2n2222

R5 output 0 10Meg


**
** Sources
**
V1 v+ 0 dc 9
V2 input 0 sin(0 0.1 1k 0 0)


**
** Models
**
.model q2n2222 npn is=19f bf=150 vaf=100 ikf=.18
+                  ise=50p ne=2.5 br=7.5 var=6.4 ikr=12m
+                  isc=8.7p nc=1.2 rb=50 re=0.4 rc=0.4 cje=26p
+                  tf=0.5n cjc=11p tr=7n xtb=1.5 kf=0.032f af=1


**
** Commands
**
*.plot tran v(input) v(output)
*.four 1k v(output)
.tran 1u 10m 0
.end

