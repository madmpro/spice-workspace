** Minimalist Discrete Power Amplifier
** A simple minimalistic design with pretty good performance.
**
** Date: 03 Mar 2018
** Author: Nathan Campos <nathan@innoveworkshop.com>

*.include ../models/bjt/npn/BC547B.mod
*.include ../models/bjt/pnp/BC557B.mod
.include ../models/tip31.mod
.include ../models/tip32.mod
.include ../models/1n4148.mod
.include ../models/bc547b.mod
.include ../models/bc557b.mod

* Input stage.
Cin input Qinb 10u
Rbias bias Qinb 10k
Qin Qvasb Qinb Qine BC557B
R1 Qine V+ 820
R2 Qvasb 0 18k
Rfb Qine dcoutput 10k

* VAS.
Cpc bout- Qvasb 5pF
Qvas bout- Qvasb 0 BC547B

* dcoutput current source and bias diodes.
Qcs1 Qcs2b Qcs2e V+ BC557B
Rcs1 Qcs2b 0 47k
Qcs2 bout+ Qcs2b Qcs2e BC557B
Rcs2 Qcs2e V+ 680
Db1 bout+ n001 1N4148
Db2 n001 bout- 1N4148

* dcoutput positive side.
Qdr1 Qoutpb bout+ dcoutput BC547B
Rdr1 Qoutpb V+ 680
Qoutp dcoutput Qoutpb V+ TIP32

* dcoutput negative side.
Qdr2 Qoutnb bout- dcoutput BC557B
Rdr2 Qoutnb 0 680
Qoutn dcoutput Qoutnb 0 TIP31

* dcoutput.
Cout dcoutput output 4700uF
Rload output 0 8

* Sources.
V1 V+ 0 dc 30V
Vin input 0 ac sin(0 1000mV 1k 0 0)
Vbias bias 0 dc 28.3V

**
** Commands
**
*.plot v(input) v(dcoutput)
*.four 1k v(dcoutput)
.tran 1u 10m 0

.end
